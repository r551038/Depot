actuateserver1
actuateserver2
