publisherpr01
publisherpr02
