server1forfiledelivery
server2forfiledelivery
server3forfiledelivery