Dbserver1
Dbserver2