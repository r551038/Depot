serverabc
serverdf
server34a
