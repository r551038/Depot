MQserver1
MQserver2
