SchedulerEnginenyp2.ny.ssmb.com
SchedulerEnginenjp2.nj.ssmb.com