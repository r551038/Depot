fonsrvnjp2
fonclnyp2
