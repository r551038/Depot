sefvertg2a.uat.mycompany.net
sefvertg2b.uat.mycompany.net
