filernjp1
filernjp2
filernyp1
filernyp2