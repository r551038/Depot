tcapplication1.eur.nsroot.net
tcapplication2.eur.nsroot.net
tcapplication32.eur.nsroot.net