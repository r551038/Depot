ServerBaseServices1
ServerBaseServices2
ServerBaseServices3
ServerBaseServices4

