CDLwebsrv1
CDLwebsrv2
CDLwebsrv3
CDwebsrva
