cnasappp1
cnasappp2
cnasappp3
cnagappp1
cnabappp1
cnwsappp1
cnwsappp2
ebasappp1
ebasappp2
ebabappp1
ebwsappp1
ebwsappp2
